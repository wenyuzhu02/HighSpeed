/home/ecelrc/students/wzhu1/HighSpeed/apr/Nov28run1_8/gscl45nm.lef