/home/ecelrc/students/wzhu1/HighSpeed/apr/Nov28run1_16/gscl45nm.lef