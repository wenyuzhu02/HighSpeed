/home/ecelrc/students/wzhu1/HighSpeed/apr/Nov28run1_4/gscl45nm.lef